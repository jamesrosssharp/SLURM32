/*
 *	multiplier placeholder
 *
 *
 */

module mult (
	input signed [31:0] A,
	input signed [31:0] B,
	output signed [63:0] out
);

assign out = A*B;

endmodule
