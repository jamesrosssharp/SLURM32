/*
 *	multiplier placeholder
 *
 *
 */

module mult (
	input signed [15:0] A,
	input signed [15:0] B,
	output signed [31:0] out
);

assign out = A*B;

endmodule
