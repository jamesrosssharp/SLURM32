/*
 *	multiplier placeholder
 *
 *
 */

module unsigned_mult (
	input [31:0] A,
	input [31:0] B,
	output [63:0] out
);

assign out = A*B;

endmodule
